** Profile: "SCHEMATIC1-opampSim"  [ C:\Users\Napoleon\Desktop\opamp\telestikos-PSpiceFiles\SCHEMATIC1\opampSim.sim ] 

** Creating circuit file "opampSim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../telestikos-pspicefiles/telestikos.lib" 
* From [PSPICE NETLIST] section of C:\Users\Napoleon\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 10 1 100meg
.TEMP 0 10 20 30 40 50 60 70
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
